// module AND(input A[0:7], input B[0:7]);
//   output out;
//   and(A[0], B[0], out);
// endmodule