module adder;

endmodule

module sub;

endmodule